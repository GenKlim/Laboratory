`timescale 1ns / 1ps

module Top(
    input BTNC,
    input BTNR,
    input CLK,
    output [6:0] SW,
    output [2:0] AN,
    output LED0
    );


endmodule
