
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity LR1_BEH is
    Port ( X : in  STD_LOGIC_VECTOR (3 downto 0);
           Y : out  STD_LOGIC_VECTOR (3 downto 0));
end LR1_BEH;

architecture Behavioral of LR1_BEH is

begin


end Behavioral;

