// Verilog test fixture created from schematic C:\Users\admin\Documents\Laboratory\Xilinxs\TA_LR_1\Main.sch - Fri May 26 20:33:45 2017

`timescale 1ns / 1ps

module Main_Main_sch_tb();

// Inputs

// Output

// Bidirs

// Instantiate the UUT
   Main UUT (
		
   );
// Initialize Inputs
   `ifdef auto_init
       initial begin
   `endif
endmodule
